package vpu_stimulus_pkg;

import uvm_pkg::*;

// Packet Sequence
`include "packet.sv"
`include "packet_sequence.sv"

endpackage
