package vpu_test_pkg;

import uvm_pkg::*;
import vpu_stimulus_pkg::*;
import vpu_env_pkg::*;

`include "test_collection.sv"

endpackage
