`include "VPU_PKG.svh"
module VPU_TOP
#(

)
(

);
    import VPU_PKG::*;
endmodule