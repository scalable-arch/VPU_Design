package vpu_env_pkg;

import uvm_pkg::*;
import vpu_stimulus_pkg::*;

`include "driver.sv"
`include "Monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "environment.sv"

endpackage
