package vpu_env_pkg;

import uvm_pkg::*;
import vpu_stimulus_pkg::*;

`include "driver.sv"
`include "input_agent.sv"
`include "reset_agent.sv"
`include "router_env.sv"

endpackage
