`include "VPU_PKG.svh"

module VPU_LANE
#(

)
(
    input   wire                            clk,
    input   wire                            rst_n,
);
    import VPU_PKG::*;
    
    
endmodule